`include "mycpu.h"
module cpu_core(
    input         clk,
    input         resetn,
    // inst sram interface
    output        inst_sram_req,
    output [ 3:0] inst_sram_wstrb,
    output [31:0] inst_sram_addr,
    output [31:0] inst_sram_wdata,
    input  [31:0] inst_sram_rdata,
    output [ 1:0] inst_sram_size,
    input         inst_sram_addr_ok,
    input         inst_sram_data_ok,
    output        inst_sram_wr,
    // data sram interface
    output        data_sram_req,
    output [ 3:0] data_sram_wstrb,
    output [31:0] data_sram_addr,
    output [31:0] data_sram_wdata,
    input  [31:0] data_sram_rdata,
    output [ 1:0] data_sram_size,
    input         data_sram_addr_ok,
    input         data_sram_data_ok,
    output        data_sram_wr,
    // trace debug interface
    output [31:0] debug_wb_pc,
    output [ 3:0] debug_wb_rf_wen,
    output [ 4:0] debug_wb_rf_wnum,
    output [31:0] debug_wb_rf_wdata
);

reg         reset;
always @(posedge clk) reset <= ~resetn; 

wire                         ds_allowin;
wire                         es_allowin;
wire                         ms_allowin;
wire                         ws_allowin;
wire                         fs_to_ds_valid;
wire                         ds_to_es_valid;
wire                         es_to_ms_valid;
wire                         ms_to_ws_valid;
wire [`FS_TO_DS_BUS_WD -1:0] fs_to_ds_bus;
wire [`DS_TO_ES_BUS_WD -1:0] ds_to_es_bus;
wire [`ES_TO_MS_BUS_WD -1:0] es_to_ms_bus;
wire [`MS_TO_WS_BUS_WD -1:0] ms_to_ws_bus;
wire [`WS_TO_RF_BUS_WD -1:0] ws_to_rf_bus;
wire [`BR_BUS_WD       -1:0] br_bus;
wire [`ES_FORWARD_WD   -1:0] es_forward;
wire [`MS_FORWARD_WD   -1:0] ms_forward;
wire [`WS_FORWARD_WD   -1:0] ws_forward;
wire                         final_ex;
wire [66                 :0] ws_to_fs_bus;
wire                         back_ertn_flush;
wire                         back_ex;
wire [63                 :0] counter;
wire                         ms_ertn_flush;
wire                         ms_to_es_valid;
wire                         ms_to_es_ex;
wire                         es_ex_detected_to_fs;

// IF stage
if_stage if_stage(
    .clk            (clk            ),
    .reset          (reset          ),
    //allowin
    .ds_allowin     (ds_allowin     ),
    //brbus
    .br_bus         (br_bus         ),
    //outputs
    .fs_to_ds_valid (fs_to_ds_valid ),
    .fs_to_ds_bus   (fs_to_ds_bus   ),
    // inst sram interface
    .inst_sram_req   (inst_sram_req   ),
    .inst_sram_wstrb  (inst_sram_wstrb  ),
    .inst_sram_addr (inst_sram_addr ),
    .inst_sram_wdata(inst_sram_wdata),
    .inst_sram_rdata(inst_sram_rdata),
    .ws_to_fs_bus   (ws_to_fs_bus   ),
    .es_forward     (es_forward     ),
    .ms_forward     (ms_forward     ),
    .ws_forward     (ws_forward     ),
    .back_ertn_flush(back_ertn_flush),
    .back_ex        (back_ex        ),
    .inst_sram_size (inst_sram_size ),
    .inst_sram_addr_ok(inst_sram_addr_ok),
    .inst_sram_data_ok(inst_sram_data_ok),
    .inst_sram_wr   (inst_sram_wr   ),
    .es_ex_detected_to_fs(es_ex_detected_to_fs)
);
// ID stage
id_stage id_stage(
    .clk            (clk            ),
    .reset          (reset          ),
    //allowin
    .es_allowin     (es_allowin     ),
    .ds_allowin     (ds_allowin     ),
    //from fs
    .fs_to_ds_valid (fs_to_ds_valid ),
    .fs_to_ds_bus   (fs_to_ds_bus   ),
    //to es
    .ds_to_es_valid (ds_to_es_valid ),
    .ds_to_es_bus   (ds_to_es_bus   ),
    //to fs
    .br_bus         (br_bus         ),
 
    //to rf: for write back
    .ws_to_rf_bus   (ws_to_rf_bus   ),
    .es_forward     (es_forward     ),
    .ms_forward     (ms_forward     ),
    .ws_forward     (ws_forward     ),
    .back_ertn_flush(back_ertn_flush),
    .back_ex        (back_ex        )
);
// EXE stage
exe_stage exe_stage(
    .clk            (clk            ),
    .reset          (reset          ),
    .final_ex       (final_ex       ),
    //allowin
    .ms_allowin     (ms_allowin     ),
    .es_allowin     (es_allowin     ),
    //from ds
    .ds_to_es_valid (ds_to_es_valid ),
    .ds_to_es_bus   (ds_to_es_bus   ),
    //to ms
    .es_to_ms_valid (es_to_ms_valid ),
    .es_to_ms_bus   (es_to_ms_bus   ),
    // data sram interface
    .data_sram_req  (data_sram_req   ),
    .data_sram_wstrb(data_sram_wstrb  ),
    .data_sram_addr (data_sram_addr ),
    .data_sram_wdata(data_sram_wdata),
    .es_forward     (es_forward     ),
    .ms_ertn_flush  (ms_ertn_flush  ),
    .ms_to_es_valid (ms_to_es_valid ),
    // counter from ws
    .es_counter     (counter        ),
    .back_ertn_flush(back_ertn_flush),
    .back_ex        (back_ex        ),
    .data_sram_size (data_sram_size ),
    .data_sram_addr_ok(data_sram_addr_ok),
    .data_sram_wr   (data_sram_wr   ),
    .ms_to_es_ex    (ms_to_es_ex    ),
    .es_ex_detected_to_fs(es_ex_detected_to_fs)
);
// MEM stage
mem_stage mem_stage(
    .clk            (clk            ),
    .reset          (reset          ),
    .final_ex       (final_ex       ),
    //allowin
    .ws_allowin     (ws_allowin     ),
    .ms_allowin     (ms_allowin     ),
    //from es
    .es_to_ms_valid (es_to_ms_valid ),
    .es_to_ms_bus   (es_to_ms_bus   ),
    //to ws
    .ms_to_ws_valid (ms_to_ws_valid ),
    .ms_to_ws_bus   (ms_to_ws_bus   ),
    //from data-sram
    .data_sram_rdata(data_sram_rdata),
    .data_sram_data_ok(data_sram_data_ok),
    .ms_forward     (ms_forward     ),
    .back_ertn_flush(back_ertn_flush),
    .ms_ertn_flush  (ms_ertn_flush  ),
    .ms_to_es_valid (ms_to_es_valid ),
    .back_ex        (back_ex        ),
    .ms_to_es_ex    (ms_to_es_ex    )
);
// WB stage
wb_stage wb_stage(
    .clk            (clk            ),
    .reset          (reset          ),
    //allowin
    .ws_allowin     (ws_allowin     ),
    //from ms
    .ms_to_ws_valid (ms_to_ws_valid ),
    .ms_to_ws_bus   (ms_to_ws_bus   ),
    .final_ex       (final_ex       ),
    //to rf: for write back
    .ws_to_rf_bus   (ws_to_rf_bus   ),
    //trace debug interface
    .debug_wb_pc      (debug_wb_pc      ),
    .debug_wb_rf_wen  (debug_wb_rf_wen  ),
    .debug_wb_rf_wnum (debug_wb_rf_wnum ),
    .debug_wb_rf_wdata(debug_wb_rf_wdata),
    .ws_forward       (ws_forward       ),
    .ws_to_fs_bus     (ws_to_fs_bus     ),
    //counter
    .counter          (counter          ),
    .back_ertn_flush  (back_ertn_flush  ),
    .back_ex          (back_ex          )
);

endmodule
